// COMMENT
// Modules
module myModule

// Imports
import v.vmod
import v.mod { a, b, c }

// Variable declarations
myVar := "Some string"
mut myVar := 12.2

// Variable assings
myVar = [1,2,3]
myVar = "a"